module moduleName (
    ports
);
    
/* wires and reg
.
.
.
 */
// from the inputs, check for the same writing location, then produce stall. and then instantiate all the modules. 
endmodule